

`ifndef BASE_PKG_SV
`define BASE_PKG_SV

package base_pkg;

   `include "base.svh"

endpackage

`endif

