library verilog;
use verilog.vl_types.all;
entity bc6502_tb is
end bc6502_tb;
