

`ifndef CPU_DUV_TOP_SV
`define CPU_DUV_TOP_SV

module cpu_duv_top(cpu_duv_if.cpu intf);

endmodule

`endif

