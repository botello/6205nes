

`ifndef TB_SVH
`define TB_SVH

   import tb_pkg::*;

   `include "base.svh"

   `include "request_item.sv"
   `include "response_item.sv"

   `include "tb_driver.sv"
   `include "tb_monitor.sv"
   `include "tb_generator.sv"
   `include "tb_scoreboard.sv"
   `include "tb_env.sv"

`endif

