

`ifndef BASE_SVH
`define BASE_SVH

   `include "object_base.sv"
   `include "component_base.sv"
   `include "item_base.sv"

`endif

