

`ifndef TB_PKG
`define TB_PKG

package tb_pkg;

   typedef logic [ 7:0] t_data;
   typedef logic [15:0] t_addr;

endpackage

`endif

