library verilog;
use verilog.vl_types.all;
entity sequencer is
    port(
        reset           : in     vl_logic;
        creset          : in     vl_logic;
        clk             : in     vl_logic;
        rdy             : in     vl_logic;
        any_int         : in     vl_logic;
        grp0            : in     vl_logic;
        grp1            : in     vl_logic;
        grp2x           : in     vl_logic;
        grp2m           : in     vl_logic;
        brk             : in     vl_logic;
        mop             : in     vl_logic;
        rti             : in     vl_logic;
        rts             : in     vl_logic;
        pul             : in     vl_logic;
        psh             : in     vl_logic;
        jsr             : in     vl_logic;
        jmp             : in     vl_logic;
        jmpi            : in     vl_logic;
        branch          : in     vl_logic;
        staxy           : in     vl_logic;
        ix              : in     vl_logic;
        iy              : in     vl_logic;
        absxy           : in     vl_logic;
        imm             : in     vl_logic;
        zpxy            : in     vl_logic;
        s_reset         : out    vl_logic;
        s_reset1        : out    vl_logic;
        s_reset2        : out    vl_logic;
        s_reset3        : out    vl_logic;
        s_nmi1          : out    vl_logic;
        s_nmi2          : out    vl_logic;
        s_nmi3          : out    vl_logic;
        s_nmi4          : out    vl_logic;
        s_nmi5          : out    vl_logic;
        s_ld_pch        : out    vl_logic;
        s_exec          : out    vl_logic;
        s_branch        : out    vl_logic;
        s_dataFetch     : out    vl_logic;
        s_update        : out    vl_logic;
        s_afterWrite    : out    vl_logic;
        s_ix1           : out    vl_logic;
        s_ix2           : out    vl_logic;
        s_iy1           : out    vl_logic;
        s_iy2           : out    vl_logic;
        s_abs1          : out    vl_logic;
        s_jmpi1         : out    vl_logic;
        s_jsr1          : out    vl_logic;
        s_jsr2          : out    vl_logic;
        s_pul           : out    vl_logic;
        s_rts1          : out    vl_logic;
        s_rts2          : out    vl_logic;
        s_rts3          : out    vl_logic;
        s_rti1          : out    vl_logic;
        s_rti2          : out    vl_logic;
        s_rti3          : out    vl_logic;
        s_sync          : out    vl_logic
    );
end sequencer;
