

`ifndef TB_PKG_SV
`define TB_PKG_SV

package tb_pkg;

   typedef logic [ 7:0] t_data;
   typedef logic [15:0] t_addr;

endpackage

`endif

